magic
tech sky130B
magscale 1 2
timestamp 1712740385
<< locali >>
rect -2070 8300 3390 8590
rect -2060 8170 -320 8300
rect -2060 4580 -780 8170
rect 1700 7990 3390 8300
rect 560 5316 782 5372
rect 2100 4570 3390 7990
rect -580 4410 -575 4460
rect 2334 4262 2344 4312
rect -2440 3940 -2250 4170
rect -330 4010 -140 4180
rect 1460 3960 1650 4170
rect 3570 3990 3760 4170
rect 1952 2078 2142 2090
rect 1952 2014 1996 2078
rect 2068 2014 2142 2078
rect -4200 1400 -1610 1430
rect -4250 20 -1610 1400
rect -1160 110 -200 250
rect 190 120 1150 260
rect 1540 100 2500 230
rect -1330 30 2670 100
rect 3240 30 5580 1390
rect -1330 20 5580 30
rect -4250 -180 5580 20
<< viali >>
rect -30 5318 14 5362
rect 1388 5312 1452 5376
rect -840 4410 -790 4460
rect -575 4410 -525 4460
rect 1861 4416 1899 4454
rect 2344 4255 2416 4327
rect 1938 3206 2158 3426
rect -832 2850 -612 3070
rect -832 1986 -612 2206
rect 1996 2006 2068 2078
<< metal1 >>
rect 1382 5382 1458 5388
rect 1382 5376 1394 5382
rect -36 5368 20 5374
rect -36 5306 20 5312
rect 1382 5312 1388 5376
rect 1382 5306 1394 5312
rect 1458 5306 1464 5382
rect 1382 5300 1458 5306
rect -846 4460 -784 4472
rect -846 4410 -840 4460
rect -790 4410 -784 4460
rect -846 4398 -784 4410
rect -581 4460 -519 4472
rect 1740 4460 1820 5940
rect -581 4410 -575 4460
rect -525 4454 1911 4460
rect -525 4416 1861 4454
rect 1899 4416 1911 4454
rect -525 4410 1911 4416
rect -581 4398 -519 4410
rect -840 4105 -790 4398
rect 2332 4327 2428 4333
rect 2332 4321 2344 4327
rect 2416 4321 2428 4327
rect 2332 4249 2338 4321
rect 2422 4249 2428 4321
rect 2338 4243 2422 4249
rect 618 4105 682 4108
rect -840 4102 682 4105
rect -840 4055 618 4102
rect 618 4032 682 4038
rect -838 3076 -606 3082
rect -838 3070 -826 3076
rect -838 2850 -832 3070
rect -838 2844 -826 2850
rect -606 2844 -600 3076
rect -838 2838 -606 2844
rect -838 2206 -606 2218
rect -838 1986 -832 2206
rect -612 1986 -606 2206
rect -838 1974 -606 1986
rect -832 960 -612 1974
rect 625 955 675 4032
rect 1932 3426 2164 3438
rect 1578 3206 1938 3426
rect 2158 3206 2164 3426
rect 1578 1864 1798 3206
rect 1932 3194 2164 3206
rect 1990 2084 2074 2090
rect 1984 2000 1990 2084
rect 2062 2078 2074 2084
rect 2068 2006 2074 2078
rect 2062 2000 2074 2006
rect 1990 1994 2074 2000
rect 1578 1644 2156 1864
rect 1936 900 2156 1644
rect 1840 490 2180 830
rect -990 260 -370 370
rect 1710 260 2330 380
rect -990 130 2330 260
<< via1 >>
rect 1394 5376 1458 5382
rect -36 5362 20 5368
rect -36 5318 -30 5362
rect -30 5318 14 5362
rect 14 5318 20 5362
rect -36 5312 20 5318
rect 1394 5312 1452 5376
rect 1452 5312 1458 5376
rect 1394 5306 1458 5312
rect 2338 4255 2344 4321
rect 2344 4255 2416 4321
rect 2416 4255 2422 4321
rect 2338 4249 2422 4255
rect 618 4038 682 4102
rect -826 3070 -606 3076
rect -826 2850 -612 3070
rect -612 2850 -606 3070
rect -826 2844 -606 2850
rect 1990 2078 2062 2084
rect 1990 2006 1996 2078
rect 1996 2006 2068 2078
rect 1990 2000 2062 2006
<< metal2 >>
rect 1394 5382 1458 5388
rect -42 5312 -36 5368
rect 20 5312 320 5368
rect -826 3076 -606 3082
rect 264 3070 320 5312
rect 1008 5312 1394 5376
rect 1008 4102 1072 5312
rect 1394 5300 1458 5306
rect 2332 4249 2338 4321
rect 2422 4249 2428 4321
rect 612 4038 618 4102
rect 682 4038 1072 4102
rect -606 2850 324 3070
rect -826 2838 -606 2844
rect 264 2078 320 2850
rect 2344 2692 2416 4249
rect 1996 2620 2416 2692
rect 1996 2090 2068 2620
rect 1990 2084 2068 2090
rect 2062 2078 2068 2084
rect 264 2006 1990 2078
rect 2062 2000 2068 2006
rect 1990 1994 2062 2000
use CNRATR_PCH_12C1F2  CNRATR_PCH_12C1F2_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform -1 0 3666 0 -1 4693
box -184 -124 2296 613
use CNRATR_PCH_12C1F2  CNRATR_PCH_12C1F2_1
timestamp 1695852000
transform 1 0 -2346 0 1 4194
box -184 -124 2296 613
use OTA  OTA_0
timestamp 1712738273
transform 1 0 470 0 1 5100
box -920 -390 1344 3290
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1705271942
transform 1 0 -1350 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1705271942
transform 1 0 0 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1705271942
transform 1 0 1350 0 1 0
box 0 0 1340 1340
use SUNTR_RPPO2  SUNTR_RPPO2_1 ~/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1712574495
transform 0 -1 5596 1 0 1370
box 0 0 2672 4236
use SUNTR_RPPO2  SUNTR_RPPO2_2
timestamp 1712574495
transform 0 1 -4270 -1 0 4042
box 0 0 2672 4236
<< labels >>
flabel locali 560 5316 782 5372 0 FreeSans 200 0 0 0 Vtail
port 3 nsew
flabel locali -1988 8424 2960 8526 0 FreeSans 200 0 0 0 VDD_1V8
port 1 nsew
flabel locali -3778 -114 5408 -4 0 FreeSans 200 0 0 0 VSS
port 2 nsew
<< end >>
