magic
tech sky130B
timestamp 1713523187
<< end >>
