*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_05_lpe.spi
#else
.include ../../../work/xsch/CNR_GR05.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0 dc 0
VDD_1V8  VDD_1V8  0 dc 1.8 
Vthreshold  Vthreshold  0 dc 0.9 
*Vreset Vreset 0 PULSE(0 1.8 0 1n 1n 10n 100n)
VPWR_UP VPWR_UP 0 PULSE(0 1.8 10n 1n 1n 10000n 10000n)

.IC v(xdut.vout)=1.8

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi



*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
*.save ${VPORTS}
.save v(xdut.vcomp)
#endif
.save all
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 1 1 1 100n 2u 0


#ifdef Debug5
tran 10p 1n 1p
*quit
#else
tran 1n 10000n 1n
write
quit
#endif

.endc

.end