*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_05_lpe.spi
#else
.include ../../../work/xsch/CNR_GR05.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0 dc 0
VDD_1V8  VDD_1V8  0 dc 1.8
*VP VP 0 dc 1.2

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VP VN VSS VDD_1V8 CNR_GR05


*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
*.save ${VPORTS}
#endif
.save all
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 10n 1u 0


#ifdef Nosweep


foreach vtemp -40 125
  option temp=$vtemp
  tran 1n 8u 1n
  write {cicname}_$vtemp
end

#else

foreach vtemp -40 -20 0 20 40 80 125
  option temp=$vtemp
*- 32*200n = 8.4 us =>
*- 64*200n = 16.8us => +5us =22us
*-  tran 1n 22u 1n
*- 128*200n = 25.6us => +5u = 31us
  tran 1n 31u 1n
*- 256*200n = 55.2us => +5us = 61us
*  tran 1n 61u 1n
  write {cicname}_$vtemp
end

#endif

quit

.endc

.end
