magic
tech sky130B
timestamp 1713364606
<< locali >>
rect -415 1590 620 1645
rect -415 1535 -135 1590
rect 340 1540 620 1590
rect -258 1318 -255 1350
rect 464 1037 490 1046
rect -293 1032 -262 1037
rect 93 460 119 486
rect -305 107 -260 134
rect 459 108 504 135
rect -41 -85 238 -81
rect 609 -85 619 -84
rect -416 -109 619 -85
<< viali >>
rect -370 1446 -340 1476
rect 544 1445 574 1476
rect -290 1318 -258 1350
rect 477 1321 503 1347
rect -373 1176 -337 1212
rect 541 1186 577 1222
rect -290 1110 -258 1142
rect -293 1037 -260 1069
rect 462 1046 498 1082
rect -292 386 -266 412
rect 461 379 491 409
rect -215 234 -179 270
rect 92 233 127 268
rect 385 236 414 265
rect 95 105 127 137
rect 98 -51 124 -25
<< metal1 >>
rect -373 1476 -337 1482
rect -373 1446 -370 1476
rect -340 1446 -337 1476
rect -373 1218 -337 1446
rect 541 1476 577 1482
rect 541 1445 544 1476
rect 574 1445 577 1476
rect -293 1350 -255 1356
rect -293 1318 -290 1350
rect -258 1347 509 1350
rect -258 1321 477 1347
rect 503 1321 509 1347
rect -258 1318 509 1321
rect -293 1312 -255 1318
rect -376 1212 -334 1218
rect -376 1176 -373 1212
rect -337 1176 -334 1212
rect -376 1170 -334 1176
rect -290 1145 -258 1312
rect 541 1225 577 1445
rect 535 1222 583 1225
rect 535 1186 541 1222
rect 577 1186 583 1222
rect 535 1183 583 1186
rect -296 1142 -252 1145
rect -296 1110 -290 1142
rect -258 1110 -252 1142
rect -296 1107 -252 1110
rect 456 1082 504 1085
rect -299 1069 -254 1072
rect -459 1037 -293 1069
rect -260 1037 -254 1069
rect 456 1046 462 1082
rect 498 1046 672 1082
rect 456 1043 504 1046
rect -459 415 -426 1037
rect -299 1034 -254 1037
rect -459 412 -260 415
rect 636 412 672 1046
rect -459 386 -292 412
rect -266 386 -260 412
rect -459 383 -260 386
rect 455 409 672 412
rect 455 379 461 409
rect 491 379 672 409
rect 455 376 672 379
rect -218 270 -176 276
rect 89 270 130 274
rect -218 234 -215 270
rect -179 268 130 270
rect -179 234 92 268
rect -218 228 -176 234
rect 89 233 92 234
rect 127 265 420 268
rect 127 236 385 265
rect 414 236 420 265
rect 127 233 420 236
rect 89 227 130 233
rect 89 137 133 140
rect 89 105 95 137
rect 127 105 133 137
rect 89 102 133 105
rect 95 -25 127 102
rect 95 -51 98 -25
rect 124 -51 127 -25
rect 95 -57 127 -51
use CNRATR_NCH_4C1F2  CNRATR_NCH_4C1F2_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -398 -1 0 634
box -92 -62 764 306
use CNRATR_NCH_4C1F2  CNRATR_NCH_4C1F2_1
timestamp 1695852000
transform 0 1 357 -1 0 634
box -92 -62 764 306
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 -1 261 1 0 -39
box -92 -62 764 364
use CNRATR_PCH_4C1F2  CNRATR_PCH_4C1F2_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 -1 -154 1 0 822
box -92 -62 764 306
use CNRATR_PCH_4C1F2  CNRATR_PCH_4C1F2_1
timestamp 1695852000
transform 0 -1 601 1 0 822
box -92 -62 764 306
<< labels >>
flabel locali 34 1594 64 1624 0 FreeSans 200 0 0 0 VDD_1V8
port 1 nsew
flabel locali 471 118 485 128 0 FreeSans 100 0 0 0 VN
port 3 nsew
flabel locali -285 116 -271 126 0 FreeSans 100 0 0 0 VP
port 4 nsew
flabel metal1 642 719 672 749 0 FreeSans 200 0 0 0 VO
port 5 nsew
flabel locali 64 -107 139 -87 0 FreeSans 400 0 0 0 VSS
port 2 nsew
flabel locali 93 460 119 486 0 FreeSans 800 0 0 0 Vtail
port 6 nsew
<< end >>
