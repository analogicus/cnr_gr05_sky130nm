magic
tech sky130B
magscale 1 2
timestamp 1713529118
<< locali >>
rect 5014 30904 5038 30944
rect 4165 12404 4646 12490
rect 5034 12404 5573 12490
rect 4165 8822 4251 12404
rect 5487 8822 5573 12404
rect 2202 8446 7660 8822
rect 4900 6221 4998 6230
rect 4900 6135 4912 6221
rect 4900 6132 4998 6135
rect 2946 -1422 3032 89
rect 6851 -1420 6937 89
rect 2944 -2160 4476 -1964
rect 5400 -2156 6940 -1966
rect -5085 -8923 -4939 -8055
rect -5085 -9057 -5079 -8923
rect -4945 -9057 -4939 -8923
rect -5085 -9063 -4939 -9057
rect -2491 -13598 -2221 -8071
rect -669 -10124 10743 -9978
rect 3920 -10412 5994 -10124
rect 12107 -13598 12377 -7771
rect 14651 -8805 14797 -7769
rect 14651 -8939 14657 -8805
rect 14791 -8939 14797 -8805
rect 14651 -8945 14797 -8939
rect -2491 -13868 4196 -13598
rect 5724 -13868 12377 -13598
<< viali >>
rect 4680 11524 4724 11568
rect 4912 6135 4998 6221
rect 1977 4357 2155 4535
rect 7681 4369 7859 4547
rect 3118 -260 3308 -70
rect 6576 -260 6766 -70
rect -5079 -9057 -4945 -8923
rect -815 -10124 -669 -9978
rect 10743 -10124 10889 -9978
rect 5678 -10849 5737 -10790
rect 4912 -11549 4998 -11463
rect 14657 -8939 14791 -8805
<< metal1 >>
rect 4674 11574 4730 11580
rect 4668 11518 4674 11574
rect 4730 11518 4736 11574
rect 4674 11512 4730 11518
rect 4806 11035 5347 11106
rect 5276 9350 5347 11035
rect 5276 9279 6281 9350
rect 4906 6227 5004 6233
rect 4900 6129 4906 6227
rect 5004 6129 5010 6227
rect 4906 6123 5004 6129
rect 1971 4535 2161 4547
rect 1971 4357 1977 4535
rect 2155 4357 2161 4535
rect 1971 -70 2161 4357
rect 6210 3790 6281 9279
rect 5947 3719 6281 3790
rect 7675 4547 7865 4559
rect 7675 4369 7681 4547
rect 7859 4369 7865 4547
rect 5947 2910 6018 3719
rect 5947 2839 7339 2910
rect 7268 524 7339 2839
rect 7268 447 7339 453
rect 3112 -70 3314 -58
rect 1971 -260 3118 -70
rect 3308 -260 3314 -70
rect 3112 -272 3314 -260
rect 6570 -70 6772 -58
rect 7675 -70 7865 4369
rect 6570 -260 6576 -70
rect 6766 -260 7865 -70
rect 6570 -272 6772 -260
rect 4906 -1556 5004 -1550
rect 4896 -1654 4906 -1558
rect 4906 -1660 5004 -1654
rect 14645 -8805 14803 -8799
rect -5091 -8923 -4933 -8917
rect -5091 -9057 -5079 -8923
rect -4945 -9057 -4933 -8923
rect 14645 -8939 14657 -8805
rect 14791 -8939 14803 -8805
rect 14645 -8945 14803 -8939
rect -5091 -9063 -4933 -9057
rect -5085 -9978 -4939 -9063
rect -821 -9978 -663 -9966
rect -5085 -10124 -815 -9978
rect -669 -10124 -663 -9978
rect -821 -10136 -663 -10124
rect 10737 -9978 10895 -9966
rect 14651 -9978 14797 -8945
rect 10737 -10124 10743 -9978
rect 10889 -10124 14797 -9978
rect 10737 -10136 10895 -10124
rect 5672 -10784 5743 -10778
rect 5666 -10855 5672 -10784
rect 5743 -10855 5749 -10784
rect 5672 -10861 5743 -10855
rect 4900 -11555 4906 -11457
rect 5004 -11555 5010 -11457
rect -2054 -12000 -1982 -11994
rect -1982 -12072 3892 -12000
rect -2054 -12078 -1982 -12072
<< via1 >>
rect 4674 11568 4730 11574
rect 4674 11524 4680 11568
rect 4680 11524 4724 11568
rect 4724 11524 4730 11568
rect 4674 11518 4730 11524
rect 4906 6221 5004 6227
rect 4906 6135 4912 6221
rect 4912 6135 4998 6221
rect 4998 6135 5004 6221
rect 4906 6129 5004 6135
rect 7268 453 7339 524
rect 4906 -1654 5004 -1556
rect 5672 -10790 5743 -10784
rect 5672 -10849 5678 -10790
rect 5678 -10849 5737 -10790
rect 5737 -10849 5743 -10790
rect 5672 -10855 5743 -10849
rect 4906 -11463 5004 -11457
rect 4906 -11549 4912 -11463
rect 4912 -11549 4998 -11463
rect 4998 -11549 5004 -11463
rect 4906 -11555 5004 -11549
rect -2054 -12072 -1982 -12000
<< metal2 >>
rect 4534 11518 4674 11574
rect 4730 11518 4736 11574
rect 4534 5486 4590 11518
rect 4911 6227 4999 6231
rect 4900 6129 4906 6227
rect 5004 6129 5010 6227
rect 4911 6125 4999 6129
rect 7262 453 7268 524
rect 7339 453 7345 524
rect 4906 -1556 5004 -1547
rect 4900 -1654 4906 -1556
rect 5004 -1654 5010 -1556
rect 4906 -1663 5004 -1654
rect 7268 -2296 7339 453
rect 5723 -2367 7339 -2296
rect -3782 -4014 -1982 -3942
rect -2054 -12000 -1982 -4014
rect 5723 -4986 5794 -2367
rect 5167 -5057 5794 -4986
rect 5167 -9666 5238 -5057
rect 5167 -9737 5743 -9666
rect 5672 -10784 5743 -9737
rect 5672 -10861 5743 -10855
rect 4906 -11457 5004 -11451
rect 4902 -11550 4906 -11462
rect 5004 -11550 5008 -11462
rect 4906 -11561 5004 -11555
rect -2060 -12072 -2054 -12000
rect -1982 -12072 -1976 -12000
<< via2 >>
rect 4911 6134 4999 6222
rect 4906 -1654 5004 -1556
rect 4911 -11550 4999 -11462
<< metal3 >>
rect 4906 6222 5004 6227
rect 4906 6134 4911 6222
rect 4999 6134 5004 6222
rect 4906 -1551 5004 6134
rect 4901 -1556 5009 -1551
rect 4901 -1654 4906 -1556
rect 5004 -1654 5009 -1556
rect 4901 -1659 5009 -1654
rect 4906 -11462 5004 -1659
rect 4906 -11550 4911 -11462
rect 4999 -11550 5004 -11462
rect 4906 -11555 5004 -11550
use INTEGRATOR  INTEGRATOR_0
timestamp 1713524416
transform 1 0 -19121 0 -1 15196
box -855 -17450 48662 6396
use IREF  IREF_0
timestamp 1713513383
transform 1 0 3800 0 1 -1114
box -3026 -8906 5302 1046
use OR  OR_0
timestamp 1713355520
transform 1 0 3068 0 1 -18806
box -184 -234 5668 4598
use OTA  OTA_0
timestamp 1713364606
transform -1 0 5164 0 -1 -10578
box -920 -262 1344 3290
use POSEDGE  POSEDGE_0
timestamp 1713520366
transform -1 0 -2158 0 1 5275
box -2052 -13405 6868 3116
use POSEDGE  POSEDGE_1
timestamp 1713520366
transform 1 0 12024 0 1 5481
box -2052 -13405 6868 3116
use PTAT  PTAT_0
timestamp 1713511997
transform 1 0 4270 0 1 180
box -4270 -180 5596 8590
<< labels >>
flabel locali 4604 8786 4754 8804 0 FreeSans 1600 0 0 0 VDD_1V8
port 1 nsew
flabel locali 7766 -10108 7968 -10042 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel locali 5014 30904 5038 30944 0 FreeSans 1600 0 0 0 RST
port 3 nsew
<< end >>
