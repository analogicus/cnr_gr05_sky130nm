magic
tech sky130B
magscale 1 2
timestamp 1713365206
<< locali >>
rect -2070 8300 3390 8590
rect -2060 8170 -320 8300
rect -2060 4718 -780 8170
rect 1700 7990 3390 8300
rect 784 6024 834 6062
rect 2100 4888 3390 7990
rect 2100 4730 3392 4888
rect 2100 4729 3762 4730
rect -2442 4614 -140 4718
rect 1458 4626 3762 4729
rect -2442 4580 -780 4614
rect -2442 4158 -1994 4580
rect 2100 4570 3762 4626
rect -580 4410 -575 4460
rect 2098 4412 2131 4484
rect 3314 4168 3762 4570
rect -4200 1400 -1610 1430
rect -4250 20 -1610 1400
rect -1160 110 -200 250
rect 190 120 1150 260
rect 1540 100 2500 230
rect -1330 30 2670 100
rect 3240 30 5580 1390
rect -1330 20 5580 30
rect -4250 -180 5580 20
<< viali >>
rect -30 5318 14 5362
rect 1388 5312 1452 5376
rect -840 4410 -790 4460
rect -575 4410 -525 4460
rect 1861 4416 1899 4454
rect 2131 4412 2204 4485
rect -832 3206 -612 3426
rect 1940 3212 2148 3420
rect -832 1986 -612 2206
rect 1938 1986 2158 2206
<< metal1 >>
rect 1382 5382 1458 5388
rect 1382 5376 1394 5382
rect -36 5368 20 5374
rect -36 5306 20 5312
rect 1382 5312 1388 5376
rect 1382 5306 1394 5312
rect 1458 5306 1464 5382
rect 1382 5300 1458 5306
rect -846 4460 -784 4472
rect -846 4410 -840 4460
rect -790 4410 -784 4460
rect -846 4398 -784 4410
rect -581 4460 -519 4472
rect 1740 4460 1820 5940
rect 2119 4485 2216 4491
rect 2119 4479 2131 4485
rect 2204 4479 2216 4485
rect -581 4410 -575 4460
rect -525 4454 1911 4460
rect -525 4416 1861 4454
rect 1899 4416 1911 4454
rect -525 4410 1911 4416
rect -581 4398 -519 4410
rect 2119 4406 2125 4479
rect 2210 4406 2216 4479
rect 2125 4400 2210 4406
rect -840 4105 -790 4398
rect 618 4105 682 4108
rect -840 4102 682 4105
rect -840 4055 618 4102
rect 618 4032 682 4038
rect -838 3432 -606 3438
rect -838 3426 -826 3432
rect -838 3206 -832 3426
rect -838 3200 -826 3206
rect -606 3200 -600 3432
rect -838 3194 -606 3200
rect -844 2206 -600 2212
rect -844 1986 -832 2206
rect -612 1986 -600 2206
rect -844 1980 -600 1986
rect -832 1916 -612 1980
rect -838 1696 -832 1916
rect -612 1696 -606 1916
rect -832 800 -612 1696
rect 625 955 675 4032
rect 1934 3426 2154 3432
rect 1934 3200 2154 3206
rect 1926 2206 2170 2212
rect 1926 1986 1938 2206
rect 2158 1986 2170 2206
rect 1926 1980 2170 1986
rect 1938 1922 2158 1980
rect 1936 1916 2158 1922
rect 2156 1696 2158 1916
rect 1936 1690 2158 1696
rect 1938 898 2158 1690
rect 1840 490 2180 830
rect -990 260 -370 370
rect 1710 260 2330 380
rect -990 130 2330 260
<< via1 >>
rect 1394 5376 1458 5382
rect -36 5362 20 5368
rect -36 5318 -30 5362
rect -30 5318 14 5362
rect 14 5318 20 5362
rect -36 5312 20 5318
rect 1394 5312 1452 5376
rect 1452 5312 1458 5376
rect 1394 5306 1458 5312
rect 2125 4412 2131 4479
rect 2131 4412 2204 4479
rect 2204 4412 2210 4479
rect 2125 4406 2210 4412
rect 618 4038 682 4102
rect -826 3426 -606 3432
rect -826 3206 -612 3426
rect -612 3206 -606 3426
rect -826 3200 -606 3206
rect -832 1696 -612 1916
rect 1934 3420 2154 3426
rect 1934 3212 1940 3420
rect 1940 3212 2148 3420
rect 2148 3212 2154 3420
rect 1934 3206 2154 3212
rect 1936 1696 2156 1916
<< metal2 >>
rect 1394 5382 1458 5388
rect -42 5312 -36 5368
rect 20 5312 320 5368
rect -826 3432 -606 3438
rect 264 3426 320 5312
rect 1008 5312 1394 5376
rect 1008 4102 1072 5312
rect 1394 5300 1458 5306
rect 2119 4406 2125 4479
rect 2210 4406 2216 4479
rect 612 4038 618 4102
rect 682 4038 1072 4102
rect 2131 3426 2204 4406
rect -606 3206 1934 3426
rect 2154 3206 2204 3426
rect 2131 3204 2204 3206
rect -826 3194 -606 3200
rect -832 1916 -612 1922
rect -612 1696 1936 1916
rect 2156 1696 2162 1916
rect -832 1690 -612 1696
use CNRATR_PCH_12C1F2  CNRATR_PCH_12C1F2_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform -1 0 3666 0 -1 4693
box -184 -124 2296 613
use CNRATR_PCH_12C1F2  CNRATR_PCH_12C1F2_1
timestamp 1695852000
transform 1 0 -2346 0 1 4194
box -184 -124 2296 613
use OTA  OTA_0
timestamp 1713364606
transform 1 0 470 0 1 5100
box -920 -262 1344 3290
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1705271942
transform 1 0 -1350 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1705271942
transform 1 0 0 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1705271942
transform 1 0 1350 0 1 0
box 0 0 1340 1340
use SUNTR_RPPO2  SUNTR_RPPO2_1 ~/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1712574495
transform 0 -1 5596 1 0 1370
box 0 0 2672 4236
use SUNTR_RPPO2  SUNTR_RPPO2_2
timestamp 1712574495
transform 0 1 -4270 1 0 1370
box 0 0 2672 4236
<< labels >>
flabel locali -1988 8424 2960 8526 0 FreeSans 200 0 0 0 VDD_1V8
port 1 nsew
flabel locali -3778 -114 5408 -4 0 FreeSans 200 0 0 0 VSS
port 2 nsew
flabel locali 784 6024 834 6062 0 FreeSans 800 0 0 0 Vtail
port 3 nsew
<< end >>
