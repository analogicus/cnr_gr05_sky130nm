*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_05_lpe.spi
#else
.include ../../../work/xsch/CNR_GR05.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0 dc 0
VDD_1V8  VDD_1V8  0 dc 1.8 
Vthreshold  Vthreshold  0 dc 1.3
VPWR_UP VPWR_UP 0 PULSE(0 1.8 10n 1n 1n 10000n 10000n)


VCLK VCLK 0 PULSE(0 1.8 0 1n 1n 10n 20n)
VA VA 0 PULSE(0 1.8 0 1n 1n 20n 40n)
*VB VB 0 PULSE(0 1.8 0 1n 1n 40n 80n)


.IC v(xdut.vout)=1.8

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

adut [VCLK VA VB] [VY] null vdut
.model vdut d_cosim simulation="./../verilog_include_file.so" 

* /home/trondfc/aicex/ip/cnr_gr05_sky130nm/sim/CNR_05/output_time
* /home/trondfc/aicex/ip/cnr_gr05_sky130nm/design/CNR_GR05_SKY130NM
* ../../../design/CNR_GR05_SKY130NM/verilog_include_file.so


*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
*.save ${VPORTS}
.save v(xdut.vcomp)
#endif
.save all
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 1 1 1 100n 2u 0


#ifdef Debug5
tran 10p 1n 1p
*quit
#else
tran 1n 1u 1n uic
write
quit
#endif

.endc

.end