** sch_path: /home/trondfc/aicex/ip/cnr_gr05_sky130nm/design/CNR_GR05_SKY130NM/CNR_GR05.sch
**.subckt CNR_GR05 VDD_1V8 VSS
*.ipin VDD_1V8
*.ipin VSS
x1 VDD_1V8 VSS VSS IREF
**** begin user architecture code


* ngspice commands
.include corner.spi


**** end user architecture code
**.ends

* expanding   symbol:  CNR_GR05_SKY130NM/IREF.sym # of pins=3
** sym_path: /home/trondfc/aicex/ip/cnr_gr05_sky130nm/design/CNR_GR05_SKY130NM/IREF.sym
** sch_path: /home/trondfc/aicex/ip/cnr_gr05_sky130nm/design/CNR_GR05_SKY130NM/IREF.sch
.subckt IREF VDD_1V8 I_REF VSS
*.ipin VDD_1V8
*.ipin VSS
*.opin I_REF
V1 net4 I_REF 0
x1 net2 net2 VDD_1V8 VDD_1V8 CNRATR_PCH_2C1F2
x2 net4 net2 VDD_1V8 VDD_1V8 CNRATR_PCH_2C1F2
x3 net3 net2 VDD_1V8 VDD_1V8 CNRATR_PCH_2C1F2
x4 net2 net3 net5 net1 CNRATR_NCH_4C8F0
x5 net3 net3 VSS VSS CNRATR_NCH_4C8F0
R1 net5 VSS 200k m=1
.ends


* expanding   symbol:  CNR_ATR_SKY130NM/CNRATR_PCH_2C1F2.sym # of pins=4
** sym_path: /home/trondfc/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_2C1F2.sym
** sch_path: /home/trondfc/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_2C1F2.sch
.subckt CNRATR_PCH_2C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.252 W=1.92 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  CNR_ATR_SKY130NM/CNRATR_NCH_4C8F0.sym # of pins=4
** sym_path: /home/trondfc/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C8F0.sym
** sch_path: /home/trondfc/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C8F0.sch
.subckt CNRATR_NCH_4C8F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=2.7 W=3.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
