*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_05_lpe.spi
#else
.include ../../../work/xsch/CNR_GR05.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0 dc 0
VDD_1V8  VDD_1V8  0 dc 1.8 
Vthreshold  Vthreshold  0 dc 1.3
VPWR_UP VPWR_UP 0 PULSE(0 1.8 10n 1n 1n 10000n 10000n)


VCLK VCLK 0 PULSE(0 1.8 0 1n 1n 12.5n 25n)
*VA VA 0 PULSE(0 1.8 200u 1n 1n 100n 200u)
*VB VB 0 PULSE(0 1.8 0 1n 1n 4000n 8000n)


.IC v(xdut.vout)=1.8

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

adut [VCLK VPWR_UP VB] [~D12 ~D11 ~D10 ~D9 ~D8 ~D7 ~D6 ~D5 ~D4 ~D3 ~D2 ~D1 ~D0] null vdut
*adut [clk reset_n signal_in] [~D7 ~D6 ~D5 ~D4 ~D3 ~D2 ~D1 ~D0] null vdut
*.model vdut d_cosim simulation="./../pulseDuration.so" 


*adut [VCLK VA VB] null null vdut
.model vdut d_cosim simulation="./../verilog_include_file.so" 



*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
*.save ${VPORTS}
.save v(xdut.vcomp)
.save v(d0)
.save v(d1)
.save v(d2)
.save v(d3)
.save v(d4)
.save v(d5)
.save v(d6)
.save v(d7)
.save v(d8)
.save v(d9)
.save v(d10)
.save v(d11)
.save v(d12)
.save v(xdut.vout)  
#endif
*.save all
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

option temp=27
optran 1 1 1 100n 2u 0


#ifdef Debug5
tran 10p 1n 1p
*quit
#else
tran 10n 250u 1n uic
write
quit
#endif

.endc

.end