magic
tech sky130B
magscale 1 2
timestamp 1713520366
<< pwell >>
rect 1392 -9196 1394 -9004
<< locali >>
rect 4224 3086 4624 3092
rect 4224 2698 4230 3086
rect 4618 2698 4624 3086
rect 4224 1312 4624 2698
rect -3 -370 2299 135
rect 2473 -355 4792 110
rect -3 -2172 2299 -1667
rect 2472 -2202 4792 -1668
rect -11 -3970 2291 -3465
rect 2468 -3976 4788 -3442
rect -10 -5394 2279 -5221
rect 20 -5729 2279 -5394
rect 2465 -5769 4785 -5235
rect 274 -7402 2291 -6945
rect 4683 -7220 4770 -6808
rect 4683 -7221 5478 -7220
rect 4683 -7607 5076 -7221
rect 5462 -7607 5478 -7221
rect 4683 -7620 5478 -7607
rect 270 -11984 350 -8723
rect 1306 -9024 1394 -9004
rect 4683 -9005 4770 -7620
rect 3475 -9197 4770 -9005
rect 2483 -11948 3592 -11656
rect 9 -13405 2307 -13131
rect 2483 -13176 3572 -13153
rect 4068 -13176 4803 -13153
rect 2483 -13400 4803 -13176
rect 2483 -13401 3572 -13400
rect 4068 -13401 4803 -13400
<< viali >>
rect 4230 2698 4618 3086
rect 5076 -7607 5462 -7221
<< metal1 >>
rect 4224 3092 4624 3098
rect 4218 2692 4224 3092
rect 4624 2692 4630 3092
rect 4224 2686 4624 2692
rect 2354 1021 2360 1052
rect 2282 985 2360 1021
rect 2427 1021 2433 1052
rect 2427 985 2509 1021
rect 2282 914 2509 985
rect -1280 -1084 -1274 -684
rect -874 -836 -868 -684
rect 2339 -773 2413 786
rect -874 -908 1060 -836
rect 5786 -842 5792 -684
rect -874 -1084 -868 -908
rect 988 -980 1060 -908
rect 3738 -914 5792 -842
rect 3738 -980 3810 -914
rect 988 -1052 1372 -980
rect 3396 -1052 3814 -980
rect -1382 -2508 -982 -2502
rect 2342 -2553 2416 -1052
rect 5786 -1084 5792 -914
rect 6192 -1084 6198 -684
rect 5814 -2478 6214 -2472
rect -982 -2720 854 -2648
rect 782 -2776 854 -2720
rect 4034 -2728 5814 -2656
rect 4034 -2776 4106 -2728
rect 782 -2848 1366 -2776
rect 2216 -2848 4106 -2776
rect -1382 -2914 -982 -2908
rect 2329 -4350 2403 -2848
rect 5814 -2884 6214 -2878
rect 2326 -6133 2403 -4571
rect 2332 -6409 2338 -6345
rect 2402 -6409 2408 -6345
rect 5070 -7215 5468 -7209
rect 5064 -7613 5070 -7215
rect 5468 -7613 5474 -7215
rect 5070 -7619 5468 -7613
rect 2427 -9279 2491 -9273
rect 2427 -9349 2491 -9343
rect 2381 -12258 2445 -12252
rect 2381 -12328 2445 -12322
rect 2262 -12718 2521 -12534
<< via1 >>
rect 4224 3086 4624 3092
rect 4224 2698 4230 3086
rect 4230 2698 4618 3086
rect 4618 2698 4624 3086
rect 4224 2692 4624 2698
rect 2360 985 2427 1052
rect -1274 -1084 -874 -684
rect -1382 -2908 -982 -2508
rect 5792 -1084 6192 -684
rect 5814 -2878 6214 -2478
rect 2338 -6409 2402 -6345
rect 5070 -7221 5468 -7215
rect 5070 -7607 5076 -7221
rect 5076 -7607 5462 -7221
rect 5462 -7607 5468 -7221
rect 5070 -7613 5468 -7607
rect 2427 -9343 2491 -9279
rect 2381 -12322 2445 -12258
<< metal2 >>
rect 4224 3092 4624 3098
rect 4220 2697 4224 3087
rect 4624 2697 4628 3087
rect 4224 2686 4624 2692
rect 2360 1109 3350 1176
rect 2360 1052 2427 1109
rect 2360 979 2427 985
rect -1274 -684 -874 -678
rect -1283 -1084 -1274 -684
rect -874 -1084 -865 -684
rect -1274 -1090 -874 -1084
rect -1382 -2508 -982 -2499
rect -1388 -2908 -1382 -2508
rect -982 -2908 -976 -2508
rect -1382 -2917 -982 -2908
rect 2338 -6345 2402 -6339
rect 2338 -6747 2402 -6409
rect 1560 -6811 2402 -6747
rect 1560 -8036 1624 -6811
rect 3283 -8001 3350 1109
rect 5792 -684 6192 -678
rect 5783 -1084 5792 -684
rect 6192 -1084 6201 -684
rect 5792 -1090 6192 -1084
rect 5814 -2478 6214 -2469
rect 5808 -2878 5814 -2478
rect 6214 -2878 6220 -2478
rect 5814 -2887 6214 -2878
rect 5075 -7215 5463 -7211
rect 5064 -7613 5070 -7215
rect 5468 -7613 5474 -7215
rect 5075 -7617 5463 -7613
rect 2204 -9343 2427 -9279
rect 2491 -9343 2497 -9279
rect 2204 -11751 2268 -9343
rect 2204 -11815 2445 -11751
rect 2381 -12258 2445 -11815
rect 2375 -12322 2381 -12258
rect 2445 -12322 2451 -12258
<< via2 >>
rect 4229 2697 4619 3087
rect -1274 -1084 -874 -684
rect -1382 -2908 -982 -2508
rect 5792 -1084 6192 -684
rect 5814 -2878 6214 -2478
rect 5075 -7608 5463 -7220
<< metal3 >>
rect 4224 3091 4624 3092
rect 4219 2693 4225 3091
rect 4623 2693 4629 3091
rect 4224 2692 4624 2693
rect -1285 -1089 -1279 -679
rect -879 -684 -869 -679
rect -874 -1084 -869 -684
rect -879 -1089 -869 -1084
rect 5787 -684 5797 -679
rect 5787 -1084 5792 -684
rect 5787 -1089 5797 -1084
rect 6197 -1089 6203 -679
rect 5809 -2478 6219 -2473
rect 5809 -2483 5814 -2478
rect 6214 -2483 6219 -2478
rect -1387 -2508 -977 -2503
rect -1387 -2513 -1382 -2508
rect -982 -2513 -977 -2508
rect 5809 -2889 6219 -2883
rect -1387 -2919 -977 -2913
rect 5071 -7215 5467 -7210
rect 5070 -7216 5468 -7215
rect 5070 -7612 5071 -7216
rect 5467 -7612 5468 -7216
rect 5070 -7613 5468 -7612
rect 5071 -7618 5467 -7613
<< via3 >>
rect 4225 3087 4623 3091
rect 4225 2697 4229 3087
rect 4229 2697 4619 3087
rect 4619 2697 4623 3087
rect 4225 2693 4623 2697
rect -1279 -684 -879 -679
rect -1279 -1084 -1274 -684
rect -1274 -1084 -879 -684
rect -1279 -1089 -879 -1084
rect 5797 -684 6197 -679
rect 5797 -1084 6192 -684
rect 6192 -1084 6197 -684
rect 5797 -1089 6197 -1084
rect -1387 -2908 -1382 -2513
rect -1382 -2908 -982 -2513
rect -982 -2908 -977 -2513
rect 5809 -2878 5814 -2483
rect 5814 -2878 6214 -2483
rect 6214 -2878 6219 -2483
rect 5809 -2883 6219 -2878
rect -1387 -2913 -977 -2908
rect 5071 -7220 5467 -7216
rect 5071 -7608 5075 -7220
rect 5075 -7608 5463 -7220
rect 5463 -7608 5467 -7220
rect 5071 -7612 5467 -7608
<< metal4 >>
rect 4224 3091 4624 3092
rect 4224 2693 4225 3091
rect 4623 2693 4624 3091
rect 4224 2692 4624 2693
rect -880 -679 -878 -678
rect -879 -1089 -878 -679
rect -880 -1090 -878 -1089
rect 5796 -679 5798 -678
rect 5796 -1089 5797 -679
rect 5796 -1090 5798 -1089
rect 5808 -2483 6220 -2482
rect 5808 -2484 5809 -2483
rect 6219 -2484 6220 -2483
rect -1388 -2513 -976 -2512
rect -1388 -2514 -1387 -2513
rect -977 -2514 -976 -2513
rect 5070 -7216 5468 -7215
rect 5070 -7612 5071 -7216
rect 5467 -7612 5468 -7216
rect 5070 -7613 5468 -7612
<< via4 >>
rect 4248 2716 4600 3068
rect -1280 -679 -880 -678
rect -1280 -1089 -1279 -679
rect -1279 -1089 -880 -679
rect -1280 -1090 -880 -1089
rect 5798 -679 6198 -678
rect 5798 -1089 6197 -679
rect 6197 -1089 6198 -679
rect 5798 -1090 6198 -1089
rect -1388 -2913 -1387 -2514
rect -1387 -2913 -977 -2514
rect -977 -2913 -976 -2514
rect 5808 -2883 5809 -2484
rect 5809 -2883 6219 -2484
rect 6219 -2883 6220 -2484
rect 5808 -2884 6220 -2883
rect -1388 -2914 -976 -2913
rect 5094 -7589 5444 -7239
<< metal5 >>
rect -378 3112 18 3116
rect -378 3110 4624 3112
rect -378 3068 5182 3110
rect -378 2716 4248 3068
rect 4600 2716 5182 3068
rect 4222 2696 5182 2716
rect 4224 2692 5176 2696
rect -1280 -654 -880 1090
rect 5798 -654 6198 1120
rect -1304 -678 -856 -654
rect -1304 -1090 -1280 -678
rect -880 -1090 -856 -678
rect -1304 -1114 -856 -1090
rect 5774 -678 6222 -654
rect 5774 -1090 5798 -678
rect 6198 -1090 6222 -678
rect 5774 -1114 6222 -1090
rect 5784 -2484 6244 -2460
rect -1412 -2514 -952 -2490
rect -1412 -2914 -1388 -2514
rect -976 -2914 -952 -2514
rect 5784 -2884 5808 -2484
rect 6220 -2884 6244 -2484
rect 5784 -2908 6244 -2884
rect -1412 -2938 -952 -2914
rect -1382 -3836 -982 -2938
rect 5814 -3786 6214 -2908
rect -645 -6058 5468 -5660
rect 5070 -7239 5468 -6058
rect 5070 -7589 5094 -7239
rect 5444 -7589 5468 -7239
rect 5070 -7613 5468 -7589
use AND  AND_0
timestamp 1713000619
transform 1 0 2470 0 1 -8788
box -2214 -2900 2108 1480
use INV  INV_0
timestamp 1712998694
transform 0 -1 4564 1 0 -13126
box -184 -238 1340 4554
use INV  INV_1
timestamp 1712998694
transform 0 -1 4554 1 0 182
box -184 -238 1340 4554
use INV  INV_2
timestamp 1712998694
transform 0 -1 4554 1 0 -1592
box -184 -238 1340 4554
use INV  INV_3
timestamp 1712998694
transform 0 -1 4552 1 0 -3388
box -184 -238 1340 4554
use INV  INV_4
timestamp 1712998694
transform 0 -1 4542 1 0 -5164
box -184 -238 1340 4554
use INV  INV_5
timestamp 1712998694
transform 0 -1 4550 1 0 -6958
box -184 -238 1340 4554
use sky130_fd_pr__cap_mim_m3_2_2Z6F9E  sky130_fd_pr__cap_mim_m3_2_2Z6F9E_0
timestamp 1713519443
transform 1 0 -925 0 1 2033
box -849 -1081 871 1081
use sky130_fd_pr__cap_mim_m3_2_2Z6F9E  sky130_fd_pr__cap_mim_m3_2_2Z6F9E_2
timestamp 1713519443
transform -1 0 5723 0 -1 2013
box -849 -1081 871 1081
use sky130_fd_pr__cap_mim_m3_2_2Z6F9E  sky130_fd_pr__cap_mim_m3_2_2Z6F9E_3
timestamp 1713519443
transform 1 0 -1203 0 1 -4749
box -849 -1081 871 1081
use sky130_fd_pr__cap_mim_m3_2_2Z6F9E  sky130_fd_pr__cap_mim_m3_2_2Z6F9E_4
timestamp 1713519443
transform -1 0 6019 0 -1 -4725
box -849 -1081 871 1081
<< labels >>
flabel locali 2848 -13354 3075 -13247 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal1 2300 -12705 2483 -12613 0 FreeSans 800 0 0 0 O
port 7 nsew
flabel metal1 2357 922 2429 959 0 FreeSans 800 0 0 0 A
port 11 nsew
flabel locali 579 -13351 806 -13244 0 FreeSans 1600 0 0 0 VDD_1V8
port 3 nsew
<< end >>
