magic
tech sky130B
magscale 1 2
timestamp 1713008575
<< locali >>
rect -6876 2368 -6750 4862
rect -4802 4670 -3484 4864
rect -3268 776 -3164 816
<< viali >>
rect -5756 4742 -5704 4794
rect -5762 4416 -5698 4480
rect -5768 4228 -5708 4288
rect -5316 3904 -5260 3960
rect -5768 3272 -5708 3332
rect -5773 3130 -5710 3193
rect -6626 2764 -6582 2808
rect -6632 1742 -6576 1798
rect -5322 1738 -5254 1806
rect -6774 1476 -6714 1536
rect -4756 1470 -4684 1542
rect -5848 1244 -5776 1316
rect -5686 1250 -5626 1310
rect -5778 950 -5690 1038
<< metal1 >>
rect -5762 4794 -5698 4806
rect -5762 4742 -5756 4794
rect -5704 4742 -5698 4794
rect -5762 4486 -5698 4742
rect -5774 4480 -5686 4486
rect -5774 4416 -5762 4480
rect -5698 4416 -5686 4480
rect -5774 4410 -5686 4416
rect -5774 4288 -5702 4300
rect -5774 4228 -5768 4288
rect -5708 4228 -5702 4288
rect -5774 3332 -5702 4228
rect -5774 3272 -5768 3332
rect -5708 3272 -5702 3332
rect -5774 3260 -5702 3272
rect -5322 3960 -5254 3972
rect -5322 3904 -5316 3960
rect -5260 3904 -5254 3960
rect -5779 3193 -5704 3205
rect -5779 3130 -5773 3193
rect -5710 3130 -5704 3193
rect -5779 3020 -5704 3130
rect -5785 2943 -5779 3020
rect -5704 2943 -5698 3020
rect -6638 2808 -6570 2814
rect -6638 2764 -6626 2808
rect -6582 2764 -6570 2808
rect -6638 2758 -6570 2764
rect -6632 1804 -6576 2758
rect -6644 1798 -6564 1804
rect -6644 1742 -6632 1798
rect -6576 1742 -6564 1798
rect -6644 1736 -6564 1742
rect -5779 1542 -5704 2943
rect -5322 1818 -5254 3904
rect -2784 2944 -2778 3019
rect -2703 2944 -2697 3019
rect -5328 1806 -5248 1818
rect -5328 1738 -5322 1806
rect -5254 1738 -5248 1806
rect -5328 1726 -5248 1738
rect -4768 1542 -4672 1548
rect -6786 1536 -4756 1542
rect -6786 1476 -6774 1536
rect -6714 1476 -4756 1536
rect -6786 1470 -4756 1476
rect -4684 1470 -4672 1542
rect -5779 1469 -5704 1470
rect -4768 1464 -4672 1470
rect -5854 1316 -5770 1328
rect -5854 1244 -5848 1316
rect -5776 1310 -5614 1316
rect -5776 1250 -5686 1310
rect -5626 1250 -5614 1310
rect -5776 1244 -5614 1250
rect -5854 1232 -5690 1244
rect -5778 1044 -5690 1232
rect -5790 1038 -5678 1044
rect -5790 950 -5778 1038
rect -5690 950 -5678 1038
rect -5790 944 -5678 950
<< via1 >>
rect -5779 2943 -5704 3020
rect -2778 2944 -2703 3019
<< metal2 >>
rect -5779 3020 -5704 3026
rect -2778 3019 -2703 3025
rect -5704 2944 -2778 3019
rect -5779 2937 -5704 2943
rect -2778 2938 -2703 2944
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 -1 -3698 1 0 942
box -184 -124 1336 2168
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_1
timestamp 1695852000
transform 0 -1 -5726 1 0 942
box -184 -124 1336 2168
use CNRATR_PCH_2C12F0  CNRATR_PCH_2C12F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -6760 -1 0 4768
box -184 -124 1336 2168
use CNRATR_PCH_2C12F0  CNRATR_PCH_2C12F0_1
timestamp 1695852000
transform 0 1 -6760 -1 0 3616
box -184 -124 1336 2168
use INV  INV_0
timestamp 1712998694
transform 1 0 -3572 0 1 988
box -184 -238 1340 4554
<< labels >>
flabel metal1 -6622 2252 -6592 2298 0 FreeSans 400 0 0 0 B
port 5 nsew
flabel metal1 -5294 2264 -5264 2310 0 FreeSans 400 0 0 0 A
port 3 nsew
flabel locali -3268 776 -3164 816 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel locali -2918 5486 -2820 5534 0 FreeSans 800 0 0 0 VDD_1V8
port 1 nsew
flabel space -3008 3240 -2974 3308 0 FreeSans 800 0 0 0 O
port 4 nsew
<< end >>
