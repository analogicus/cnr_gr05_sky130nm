magic
tech sky130B
magscale 1 2
timestamp 1713355520
<< locali >>
rect 4236 4538 5580 4598
rect 700 3988 802 3990
rect 700 3796 918 3988
rect 2994 3796 4396 3988
rect 700 2836 802 3796
rect 700 2644 922 2836
rect 700 1684 802 2644
rect 700 1492 916 1684
rect 4036 1116 4266 1308
rect 4032 -234 4424 156
<< viali >>
rect 1956 3870 2008 3922
rect 1950 3540 2014 3604
rect 1948 3294 2000 3346
rect 1070 3028 1134 3092
rect 1942 2388 2006 2452
rect 1948 2156 2000 2208
rect 2806 1876 2870 1940
rect 1076 866 1128 918
rect 2812 868 2864 920
rect 927 542 991 610
rect 2966 550 3018 602
rect 942 348 1006 412
rect 2956 348 3020 412
rect 948 34 1000 86
rect 2962 34 3014 86
<< metal1 >>
rect 1950 3922 2014 3934
rect 1950 3870 1956 3922
rect 2008 3870 2014 3922
rect 1950 3610 2014 3870
rect 1938 3604 2026 3610
rect 1938 3540 1950 3604
rect 2014 3540 2026 3604
rect 1938 3534 2026 3540
rect 1942 3346 2006 3358
rect 1942 3294 1948 3346
rect 2000 3294 2006 3346
rect 1058 3092 1146 3098
rect 1058 3028 1070 3092
rect 1134 3028 1146 3092
rect 1058 3022 1146 3028
rect 1070 1466 1134 3022
rect 1942 2458 2006 3294
rect 1930 2452 2018 2458
rect 1930 2388 1942 2452
rect 2006 2388 2018 2452
rect 1930 2382 2018 2388
rect 1942 2208 2006 2220
rect 1942 2156 1948 2208
rect 2000 2156 2006 2208
rect 1942 1800 2006 2156
rect 4780 2020 4876 2274
rect 5134 2190 5198 2196
rect 5134 2120 5198 2126
rect 2794 1940 2882 1946
rect 2794 1876 2806 1940
rect 2870 1876 2882 1940
rect 2794 1870 2882 1876
rect 1936 1736 1942 1800
rect 2006 1736 2012 1800
rect 1070 1340 1226 1466
rect 1070 924 1134 1340
rect 1064 918 1140 924
rect 1064 866 1076 918
rect 1128 866 1140 918
rect 1064 860 1140 866
rect 921 610 997 622
rect 921 542 927 610
rect 991 608 997 610
rect 1942 608 2006 1736
rect 2806 1472 2870 1870
rect 2806 1332 2986 1472
rect 2806 920 2870 1332
rect 2806 868 2812 920
rect 2864 868 2870 920
rect 2806 856 2870 868
rect 991 602 3030 608
rect 991 550 2966 602
rect 3018 550 3030 602
rect 991 544 3030 550
rect 991 542 997 544
rect 921 530 997 542
rect 930 412 1018 418
rect 930 348 942 412
rect 1006 348 1018 412
rect 930 342 1018 348
rect 2944 412 3032 418
rect 2944 348 2956 412
rect 3020 348 3032 412
rect 2944 342 3032 348
rect 942 86 1006 342
rect 942 34 948 86
rect 1000 34 1006 86
rect 942 22 1006 34
rect 2956 86 3020 342
rect 2956 34 2962 86
rect 3014 34 3020 86
rect 2956 22 3020 34
<< via1 >>
rect 5134 2126 5198 2190
rect 1942 1736 2006 1800
<< metal2 >>
rect 3980 2126 5134 2190
rect 5198 2126 5204 2190
rect 1942 1800 2006 1806
rect 3980 1800 4044 2126
rect 2006 1736 4044 1800
rect 1942 1730 2006 1736
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 -1 4014 1 0 60
box -184 -124 1336 2168
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_1
timestamp 1695852000
transform 0 -1 1984 1 0 60
box -184 -124 1336 2168
use CNRATR_PCH_2C12F0  CNRATR_PCH_2C12F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 948 -1 0 3892
box -184 -124 1336 2168
use CNRATR_PCH_2C12F0  CNRATR_PCH_2C12F0_1
timestamp 1695852000
transform 0 1 948 -1 0 2740
box -184 -124 1336 2168
use INV  INV_0
timestamp 1712998694
transform 1 0 4328 0 1 4
box -184 -238 1340 4554
<< labels >>
flabel locali 4846 4572 4896 4586 0 FreeSans 400 0 0 0 VDD_1V8
port 1 nsew
flabel locali 4088 -162 4154 -82 0 FreeSans 400 0 0 0 VSS
port 2 nsew
flabel metal1 4800 2212 4832 2246 0 FreeSans 400 0 0 0 O
port 4 nsew
flabel metal1 2900 1366 2944 1434 0 FreeSans 400 0 0 0 B
port 5 nsew
flabel metal1 1158 1372 1200 1426 0 FreeSans 400 0 0 0 A
port 3 nsew
<< end >>
