magic
tech sky130B
timestamp 1713513383
<< locali >>
rect -340 503 1484 523
rect -340 473 271 503
rect 301 502 1484 503
rect 301 476 847 502
rect 873 476 1484 502
rect 301 473 1484 476
rect -340 462 1484 473
rect 845 424 876 426
rect 844 213 846 247
rect 269 -207 524 -111
rect 620 -207 809 -111
rect 1126 -265 1152 -262
rect 1126 -297 1152 -295
rect -19 -404 -15 -371
rect 1122 -373 1152 -369
rect 1122 -405 1152 -403
rect 245 -783 341 -422
rect 636 -436 666 -434
rect 636 -473 666 -472
rect 802 -783 898 -409
rect 245 -847 434 -783
rect 711 -847 899 -783
rect 245 -992 899 -847
rect 245 -1070 434 -992
rect 711 -1070 899 -992
rect 390 -1735 410 -1070
rect 746 -1735 766 -1070
rect 390 -1742 766 -1735
rect 409 -1831 747 -1742
rect 206 -2239 316 -1852
<< viali >>
rect 271 473 301 503
rect 847 476 873 502
rect 268 395 304 431
rect 844 392 876 424
rect 396 360 428 392
rect 719 363 745 389
rect 179 215 209 245
rect 719 215 749 245
rect 846 212 882 248
rect 1125 221 1149 245
rect 117 -256 153 -220
rect 993 -253 1023 -223
rect -91 -296 -59 -264
rect 1122 -295 1152 -265
rect 120 -346 146 -320
rect 557 -336 587 -306
rect -15 -406 21 -370
rect 1122 -403 1152 -373
rect 554 -471 590 -435
rect 633 -472 669 -436
rect 563 -1199 593 -1169
rect 560 -1332 596 -1296
rect 563 -1550 595 -1518
rect 566 -1707 592 -1681
rect 864 -2193 888 -2169
rect 206 -4118 316 -4008
rect 825 -4115 929 -4011
<< metal1 >>
rect 268 503 304 509
rect 268 473 271 503
rect 301 473 304 503
rect 268 434 304 473
rect 844 502 876 508
rect 844 476 847 502
rect 873 476 876 502
rect 262 431 310 434
rect 262 395 268 431
rect 304 395 310 431
rect 844 427 876 476
rect 838 424 882 427
rect 262 392 310 395
rect 393 392 431 398
rect 454 394 490 397
rect 393 360 396 392
rect 428 360 454 392
rect 393 354 431 360
rect 838 392 844 424
rect 876 392 882 424
rect 490 389 751 392
rect 838 389 882 392
rect 490 363 719 389
rect 745 363 751 389
rect 490 360 751 363
rect 454 355 490 358
rect 176 245 212 251
rect 843 248 885 254
rect 176 215 179 245
rect 209 215 212 245
rect 114 -220 156 -214
rect 176 -220 212 215
rect 713 245 846 248
rect 713 215 719 245
rect 749 215 846 245
rect 713 212 846 215
rect 882 212 885 248
rect 843 206 885 212
rect 1122 245 1152 251
rect 1122 221 1125 245
rect 1149 221 1152 245
rect 114 -256 117 -220
rect 153 -223 1029 -220
rect 153 -253 993 -223
rect 1023 -253 1029 -223
rect 153 -256 1029 -253
rect -97 -264 -53 -261
rect 114 -262 156 -256
rect -97 -296 -91 -264
rect -59 -296 -53 -264
rect -97 -299 -53 -296
rect -91 -317 -59 -299
rect 554 -306 590 -300
rect -91 -320 152 -317
rect -91 -346 120 -320
rect 146 -346 152 -320
rect -91 -349 152 -346
rect 554 -336 557 -306
rect 587 -336 590 -306
rect -21 -370 27 -367
rect 554 -369 590 -336
rect -21 -406 -15 -370
rect 21 -406 27 -370
rect 551 -405 554 -369
rect 590 -405 593 -369
rect -21 -409 27 -406
rect -15 -1232 21 -409
rect 554 -432 590 -405
rect 548 -435 596 -432
rect 548 -471 554 -435
rect 590 -471 596 -435
rect 548 -474 596 -471
rect 630 -436 672 -430
rect 720 -436 756 -256
rect 1122 -262 1152 221
rect 1116 -265 1158 -262
rect 1116 -295 1122 -265
rect 1152 -295 1158 -265
rect 1116 -298 1158 -295
rect 1119 -373 1155 -367
rect 1119 -403 1122 -373
rect 1152 -403 1155 -373
rect 1119 -409 1155 -403
rect 630 -472 633 -436
rect 669 -472 756 -436
rect 630 -478 672 -472
rect 560 -1169 596 -1163
rect 560 -1199 563 -1169
rect 593 -1199 596 -1169
rect 560 -1232 596 -1199
rect -15 -1268 596 -1232
rect 560 -1293 596 -1268
rect 554 -1296 602 -1293
rect 554 -1332 560 -1296
rect 596 -1332 602 -1296
rect 554 -1335 602 -1332
rect 557 -1518 601 -1515
rect 557 -1550 563 -1518
rect 595 -1550 601 -1518
rect 557 -1553 601 -1550
rect 563 -1681 595 -1553
rect 563 -1707 566 -1681
rect 592 -1707 595 -1681
rect 563 -1713 595 -1707
rect 1122 -2011 1152 -409
rect 861 -2041 1152 -2011
rect 861 -2169 891 -2041
rect 861 -2193 864 -2169
rect 888 -2193 891 -2169
rect 861 -2199 891 -2193
rect 203 -4008 319 -4002
rect 203 -4118 206 -4008
rect 316 -4011 935 -4008
rect 316 -4115 825 -4011
rect 929 -4115 935 -4011
rect 316 -4118 935 -4115
rect 203 -4124 319 -4118
<< via1 >>
rect 454 358 490 394
rect 554 -405 590 -369
<< metal2 >>
rect 451 358 454 394
rect 490 358 493 394
rect 454 -369 490 358
rect 554 -369 590 -366
rect 454 -405 554 -369
rect 554 -408 590 -405
use CNRATR_NCH_4C1F2  CNRATR_NCH_4C1F2_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 -1 694 1 0 -831
box -92 -62 764 306
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 -1 729 1 0 -1694
box -92 -62 764 364
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_1
timestamp 1695852000
transform -1 0 1522 0 -1 -128
box -92 -62 764 364
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_3
timestamp 1695852000
transform 1 0 -379 0 1 -431
box -92 -62 764 364
use CNRATR_PCH_8C4F0  CNRATR_PCH_8C4F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform -1 0 1436 0 -1 453
box -92 -62 956 508
use CNRATR_PCH_8C4F0  CNRATR_PCH_8C4F0_1
timestamp 1695852000
transform 1 0 -292 0 1 7
box -92 -62 956 508
use SUNTR_RPPO8  SUNTR_RPPO8_0 ~/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1713363649
transform 0 -1 2651 1 0 -4453
box 0 0 2632 2118
use SUNTR_RPPO8  SUNTR_RPPO8_1
timestamp 1713363649
transform 0 1 -1513 -1 0 -1821
box 0 0 2632 2118
<< labels >>
flabel metal1 559 -249 594 -232 0 FreeSans 100 0 0 0 Vref
port 3 nsew
flabel locali -214 486 -179 503 0 FreeSans 400 0 0 0 VDD_1V8
port 1 nsew
flabel locali 533 -1809 632 -1766 0 FreeSans 800 0 0 0 VSS
port 2 nsew
<< end >>
