*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/final_lpe.spi
#else
.include ../../../work/xsch/final.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0 dc 0
VDD_1V8  VDD_1V8  0 dc 1.8 
*Vthreshold  Vthreshold  0 dc 1.3
VPWR_UP VPWR_UP 0 PULSE(0 1.8 10n 1n 1n 10000n 10000n)


VCLK VCLK 0 PULSE(0 1.8 0 1n 1n 12.5n 25n)
*VA VA 0 PULSE(0 1.8 200u 1n 1n 100n 200u)
*VB VB 0 PULSE(0 1.8 0 1n 1n 4000n 8000n)


.IC v(xdut.vout)=1.8

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

adut [VCLK VPWR_UP pulse] [N] null vdut
.model vdut d_cosim simulation="./../verilog_include_file.so" 


*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
*.save ${VPORTS}
#endif
.save all
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

*option temp=-40
optran 1 1 1 100n 2u 0



tran 10n 150u 1n uic
write
quit

.endc

.end