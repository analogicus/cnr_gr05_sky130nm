magic
tech sky130B
magscale 1 2
timestamp 1713532653
<< locali >>
rect 3998 30952 4710 30958
rect 3998 30892 4004 30952
rect 4064 30892 4710 30952
rect 5014 30904 5038 30944
rect 3998 30886 4710 30892
rect 4165 12404 4646 12490
rect 5034 12404 5573 12490
rect 4165 8822 4251 12404
rect 5487 8822 5573 12404
rect 2202 8446 7660 8822
rect 4900 6221 4998 6230
rect 4900 6135 4912 6221
rect 4900 6132 4998 6135
rect -2198 5584 2352 5954
rect 7514 5782 12064 6152
rect 2946 -1422 3032 89
rect 6851 -1420 6937 89
rect 2944 -2160 4476 -1964
rect 5400 -2156 6940 -1966
rect -5085 -8923 -4939 -8055
rect -5085 -9057 -5079 -8923
rect -4945 -9057 -4939 -8923
rect -5085 -9063 -4939 -9057
rect -2491 -13598 -2221 -8071
rect -669 -10124 1884 -9978
rect 2092 -10124 10743 -9978
rect 3920 -10412 5994 -10124
rect 2424 -10714 4334 -10708
rect 2424 -10922 2430 -10714
rect 2638 -10922 4334 -10714
rect 2424 -10928 4334 -10922
rect 12107 -13598 12377 -7771
rect 14651 -8805 14797 -7769
rect 14651 -8939 14657 -8805
rect 14791 -8939 14797 -8805
rect 14651 -8945 14797 -8939
rect -2491 -13862 4235 -13598
rect 5849 -13602 12377 -13598
rect 5849 -13810 9642 -13602
rect 9850 -13810 12377 -13602
rect -2491 -13866 4456 -13862
rect 5849 -13866 12377 -13810
rect -2491 -13868 12377 -13866
rect 2972 -14254 7852 -13868
rect 4198 -14906 7852 -14254
rect 2060 -15402 2654 -15092
rect 1638 -17630 1750 -17618
rect 1586 -17724 1782 -17630
rect 1638 -19678 1750 -17724
rect 10010 -19678 10122 -17090
rect 1638 -19790 10122 -19678
<< viali >>
rect 4004 30892 4064 30952
rect 4680 11524 4724 11568
rect 4912 6135 4998 6221
rect 1977 4357 2155 4535
rect 7681 4369 7859 4547
rect 3118 -260 3308 -70
rect 6576 -260 6766 -70
rect -5079 -9057 -4945 -8923
rect -815 -10124 -669 -9978
rect 1884 -10126 2092 -9918
rect 10743 -10124 10889 -9978
rect 2430 -10922 2638 -10714
rect 5678 -10849 5737 -10790
rect 4912 -11549 4998 -11463
rect 14657 -8939 14791 -8805
rect 9642 -13810 9850 -13602
rect 1878 -15062 2098 -14842
rect 9636 -15406 9856 -15186
rect 9636 -16596 9856 -16376
rect 1896 -17110 2104 -16902
rect 8447 -18837 8581 -18703
<< metal1 >>
rect 3998 30958 4070 30964
rect 3992 30886 3998 30958
rect 4070 30886 4076 30958
rect 3998 30880 4070 30886
rect 4674 11574 4730 11580
rect 4668 11518 4674 11574
rect 4730 11518 4736 11574
rect 4674 11512 4730 11518
rect 4806 11035 5347 11106
rect 5276 9350 5347 11035
rect 5276 9279 6281 9350
rect 4906 6227 5004 6233
rect 4900 6129 4906 6227
rect 5004 6129 5010 6227
rect 4906 6123 5004 6129
rect 1971 4535 2161 4547
rect 1971 4357 1977 4535
rect 2155 4357 2161 4535
rect 1971 -70 2161 4357
rect 6210 3790 6281 9279
rect 5947 3719 6281 3790
rect 7675 4547 7865 4559
rect 7675 4369 7681 4547
rect 7859 4369 7865 4547
rect 5947 2910 6018 3719
rect 5947 2839 7339 2910
rect 7268 524 7339 2839
rect 7268 447 7339 453
rect 3112 -70 3314 -58
rect 1971 -260 3118 -70
rect 3308 -260 3314 -70
rect 3112 -272 3314 -260
rect 6570 -70 6772 -58
rect 7675 -70 7865 4369
rect 6570 -260 6576 -70
rect 6766 -260 7865 -70
rect 6570 -272 6772 -260
rect 4906 -1556 5004 -1550
rect 4896 -1654 4906 -1558
rect 4906 -1660 5004 -1654
rect 14361 -7239 14367 -7113
rect 14493 -7239 14499 -7113
rect -4636 -7452 -4630 -7312
rect -4490 -7452 -4484 -7312
rect 14645 -8805 14803 -8799
rect -5091 -8923 -4933 -8917
rect -5091 -9057 -5079 -8923
rect -4945 -9057 -4933 -8923
rect 14645 -8939 14657 -8805
rect 14791 -8939 14803 -8805
rect 14645 -8945 14803 -8939
rect -5091 -9063 -4933 -9057
rect -5085 -9978 -4939 -9063
rect 1872 -9918 2104 -9912
rect -821 -9978 -663 -9966
rect -5085 -10124 -815 -9978
rect -669 -10124 -663 -9978
rect -821 -10136 -663 -10124
rect 1872 -10126 1884 -9918
rect 2092 -10126 2104 -9918
rect 1872 -10132 2104 -10126
rect 10737 -9978 10895 -9966
rect 14651 -9978 14797 -8945
rect 10737 -10124 10743 -9978
rect 10889 -10124 14797 -9978
rect 1878 -11628 2098 -10132
rect 10737 -10136 10895 -10124
rect 2424 -10708 2644 -10702
rect 2418 -10928 2424 -10708
rect 2644 -10928 2650 -10708
rect 5672 -10784 5743 -10778
rect 5666 -10855 5672 -10784
rect 5743 -10855 5749 -10784
rect 5672 -10861 5743 -10855
rect 2424 -10934 2644 -10928
rect 4900 -11555 4906 -11457
rect 5004 -11555 5010 -11457
rect 1872 -11848 1878 -11628
rect 2098 -11848 2104 -11628
rect 1878 -11854 2098 -11848
rect -2054 -12000 -1982 -11994
rect -1982 -12072 3892 -12000
rect -2054 -12078 -1982 -12072
rect 690 -12598 696 -12378
rect 916 -12598 922 -12378
rect 1878 -12512 2098 -12506
rect 696 -17308 916 -12598
rect 1878 -14836 2098 -12732
rect 9636 -13596 9856 -13590
rect 9630 -13816 9636 -13596
rect 9856 -13816 9862 -13596
rect 9636 -13822 9856 -13816
rect 12711 -14277 12857 -10124
rect 8835 -14423 12857 -14277
rect 1866 -14842 2110 -14836
rect 1866 -15062 1878 -14842
rect 2098 -15062 2110 -14842
rect 1866 -15068 2110 -15062
rect 4868 -15584 4940 -15578
rect 3612 -15656 4868 -15584
rect 4868 -15662 4940 -15656
rect 1890 -16902 2110 -16890
rect 1890 -17110 1896 -16902
rect 2104 -17110 2110 -16902
rect 1890 -17308 2110 -17110
rect 696 -17528 2110 -17308
rect 5566 -17474 5572 -17334
rect 5712 -17474 5718 -17334
rect 7320 -17466 7326 -17340
rect 7452 -17466 7458 -17340
rect 1890 -19214 2110 -17528
rect 8835 -18697 8981 -14423
rect 9630 -15180 9862 -15174
rect 9624 -15400 9630 -15180
rect 9862 -15400 9868 -15180
rect 9624 -15406 9636 -15400
rect 9856 -15406 9868 -15400
rect 9624 -15412 9868 -15406
rect 9624 -16376 9868 -16370
rect 9624 -16596 9636 -16376
rect 9856 -16596 9868 -16376
rect 9624 -16602 9868 -16596
rect 8435 -18703 8981 -18697
rect 8435 -18837 8447 -18703
rect 8581 -18837 8981 -18703
rect 8435 -18843 8981 -18837
rect 9636 -19214 9856 -16602
rect 1890 -19434 9856 -19214
<< via1 >>
rect 3998 30952 4070 30958
rect 3998 30892 4004 30952
rect 4004 30892 4064 30952
rect 4064 30892 4070 30952
rect 3998 30886 4070 30892
rect 4674 11568 4730 11574
rect 4674 11524 4680 11568
rect 4680 11524 4724 11568
rect 4724 11524 4730 11568
rect 4674 11518 4730 11524
rect 4906 6221 5004 6227
rect 4906 6135 4912 6221
rect 4912 6135 4998 6221
rect 4998 6135 5004 6221
rect 4906 6129 5004 6135
rect 7268 453 7339 524
rect 4906 -1654 5004 -1556
rect 14367 -7239 14493 -7113
rect -4630 -7452 -4490 -7312
rect 2424 -10714 2644 -10708
rect 2424 -10922 2430 -10714
rect 2430 -10922 2638 -10714
rect 2638 -10922 2644 -10714
rect 2424 -10928 2644 -10922
rect 5672 -10790 5743 -10784
rect 5672 -10849 5678 -10790
rect 5678 -10849 5737 -10790
rect 5737 -10849 5743 -10790
rect 5672 -10855 5743 -10849
rect 4906 -11463 5004 -11457
rect 4906 -11549 4912 -11463
rect 4912 -11549 4998 -11463
rect 4998 -11549 5004 -11463
rect 4906 -11555 5004 -11549
rect 1878 -11848 2098 -11628
rect -2054 -12072 -1982 -12000
rect 696 -12598 916 -12378
rect 1878 -12732 2098 -12512
rect 9636 -13602 9856 -13596
rect 9636 -13810 9642 -13602
rect 9642 -13810 9850 -13602
rect 9850 -13810 9856 -13602
rect 9636 -13816 9856 -13810
rect 4868 -15656 4940 -15584
rect 5572 -17474 5712 -17334
rect 7326 -17466 7452 -17340
rect 9630 -15186 9862 -15180
rect 9630 -15400 9636 -15186
rect 9636 -15400 9856 -15186
rect 9856 -15400 9862 -15186
<< metal2 >>
rect 3992 30886 3998 30958
rect 4070 30886 4076 30958
rect 3998 9038 4070 30886
rect 3702 8966 4070 9038
rect 4534 11518 4674 11574
rect 4730 11518 4736 11574
rect 3702 8258 3774 8966
rect 1682 8186 3774 8258
rect 1682 1804 1754 8186
rect 4534 5486 4590 11518
rect 14362 6566 14488 6688
rect 4911 6227 4999 6231
rect 4900 6129 4906 6227
rect 5004 6129 5010 6227
rect 4911 6125 4999 6129
rect 1682 1734 2872 1804
rect 1754 1732 2872 1734
rect -5488 -972 -1982 -900
rect -4630 -7312 -4490 -7306
rect -4630 -8280 -4490 -7452
rect -4630 -8420 -2764 -8280
rect -2904 -13984 -2764 -8420
rect -2054 -12000 -1982 -972
rect 2800 -2214 2872 1732
rect 7262 453 7268 524
rect 7339 453 7345 524
rect 4906 -1556 5004 -1547
rect 4900 -1654 4906 -1556
rect 5004 -1654 5010 -1556
rect 4906 -1663 5004 -1654
rect 2800 -2286 3718 -2214
rect 1060 -10716 2424 -10708
rect 696 -10928 2424 -10716
rect 2644 -10928 2650 -10708
rect 696 -10936 1338 -10928
rect -2060 -12072 -2054 -12000
rect -1982 -12072 -1976 -12000
rect 696 -12378 916 -10936
rect 1878 -11628 2098 -11622
rect 1878 -12512 2098 -11848
rect 3646 -12348 3718 -2286
rect 7268 -2296 7339 453
rect 5723 -2367 7339 -2296
rect 5723 -4986 5794 -2367
rect 5167 -5057 5794 -4986
rect 5167 -9666 5238 -5057
rect 14367 -7113 14493 -7107
rect 14367 -8057 14493 -7239
rect 12473 -8183 14493 -8057
rect 5167 -9737 5743 -9666
rect 5672 -10784 5743 -9737
rect 5672 -10861 5743 -10855
rect 4906 -11457 5004 -11451
rect 4902 -11550 4906 -11462
rect 5004 -11550 5008 -11462
rect 4906 -11561 5004 -11555
rect 3646 -12420 4940 -12348
rect 696 -12604 916 -12598
rect 1872 -12732 1878 -12512
rect 2098 -12732 2104 -12512
rect -2904 -14124 2910 -13984
rect 2770 -17334 2910 -14124
rect 4868 -15584 4940 -12420
rect 9630 -13816 9636 -13596
rect 9856 -13816 9862 -13596
rect 12473 -13985 12599 -8183
rect 7911 -14111 12599 -13985
rect 4862 -15656 4868 -15584
rect 4940 -15656 4946 -15584
rect 5572 -17334 5712 -17328
rect 2770 -17474 5572 -17334
rect 7326 -17340 7452 -17334
rect 7911 -17340 8037 -14111
rect 9630 -15180 9862 -15171
rect 9624 -15400 9630 -15180
rect 9862 -15400 9868 -15180
rect 9630 -15409 9862 -15400
rect 7452 -17466 8037 -17340
rect 7326 -17472 7452 -17466
rect 5572 -17480 5712 -17474
<< via2 >>
rect 4911 6134 4999 6222
rect 4906 -1654 5004 -1556
rect 4911 -11550 4999 -11462
rect 9641 -13811 9851 -13601
rect 9630 -15400 9862 -15180
<< metal3 >>
rect 4906 6222 5004 6227
rect 4906 6134 4911 6222
rect 4999 6134 5004 6222
rect 4906 -1551 5004 6134
rect 4901 -1556 5009 -1551
rect 4901 -1654 4906 -1556
rect 5004 -1654 5009 -1556
rect 4901 -1659 5009 -1654
rect 4906 -11462 5004 -1659
rect 4906 -11550 4911 -11462
rect 4999 -11550 5004 -11462
rect 4906 -11555 5004 -11550
rect 9636 -13601 9856 -13596
rect 9636 -13811 9641 -13601
rect 9851 -13811 9856 -13601
rect 9636 -15175 9856 -13811
rect 9625 -15180 9867 -15175
rect 9625 -15400 9630 -15180
rect 9862 -15400 9867 -15180
rect 9625 -15405 9867 -15400
use INTEGRATOR  INTEGRATOR_0
timestamp 1713524416
transform 1 0 -19121 0 -1 15196
box -855 -17450 48662 6396
use IREF  IREF_0
timestamp 1713513383
transform 1 0 3800 0 1 -1114
box -3026 -8906 5302 1046
use OR  OR_0
timestamp 1713355520
transform -1 0 8552 0 1 -18806
box -184 -234 5668 4598
use OTA  OTA_0
timestamp 1713364606
transform -1 0 5164 0 -1 -10578
box -920 -262 1344 3290
use POSEDGE  POSEDGE_0
timestamp 1713520366
transform -1 0 -2158 0 1 5275
box -2052 -13405 6868 3116
use POSEDGE  POSEDGE_1
timestamp 1713520366
transform 1 0 12024 0 1 5481
box -2052 -13405 6868 3116
use PTAT  PTAT_0
timestamp 1713511997
transform 1 0 4270 0 1 180
box -4270 -180 5596 8590
use SUNTR_RPPO2  SUNTR_RPPO2_0 ~/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1712574495
transform 0 -1 13294 1 0 -17212
box 0 0 2672 4236
use SUNTR_RPPO4  SUNTR_RPPO4_0 ~/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1713532524
transform 0 1 -1560 -1 0 -14210
box 0 0 3536 4236
<< labels >>
flabel locali 4604 8786 4754 8804 0 FreeSans 1600 0 0 0 VDD_1V8
port 1 nsew
flabel locali 7766 -10108 7968 -10042 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal2 14408 6664 14444 6678 0 FreeSans 1600 0 0 0 VPWR_UP
port 7 nsew
<< end >>
