magic
tech sky130B
magscale 1 2
timestamp 1711874809
<< pwell >>
rect -90 -180 470 -30
<< locali >>
rect -90 2379 1220 2390
rect -90 2370 911 2379
rect -90 2310 158 2370
rect 218 2321 911 2370
rect 969 2321 1220 2379
rect 218 2310 1220 2321
rect -90 2290 1220 2310
rect -90 -170 470 -30
rect 660 -158 1220 -40
rect 660 -170 1060 -158
rect -180 -221 1060 -170
rect 1123 -170 1220 -158
rect 1123 -221 1310 -170
rect -180 -250 1310 -221
<< viali >>
rect 158 2310 218 2370
rect 911 2321 969 2379
rect 152 1660 224 1732
rect 905 1665 975 1735
rect 148 613 202 667
rect 303 608 378 683
rect 1054 614 1129 689
rect 140 327 210 393
rect 890 330 961 401
rect 1060 -221 1123 -158
<< metal1 >>
rect 152 2370 224 2382
rect 152 2310 158 2370
rect 218 2310 224 2370
rect 152 1744 224 2310
rect 905 2379 975 2391
rect 905 2321 911 2379
rect 969 2321 975 2379
rect 146 1732 230 1744
rect 905 1741 975 2321
rect 146 1660 152 1732
rect 224 1660 230 1732
rect 146 1648 230 1660
rect 893 1735 987 1741
rect 893 1665 905 1735
rect 975 1665 987 1735
rect 893 1659 987 1665
rect 297 683 384 695
rect 1042 689 1141 695
rect 1042 683 1054 689
rect 142 667 208 679
rect 142 613 148 667
rect 202 613 208 667
rect 142 525 208 613
rect 297 608 303 683
rect 378 614 1054 683
rect 1129 614 1141 689
rect 378 608 1141 614
rect 297 596 384 608
rect 135 454 961 525
rect 142 399 208 454
rect 890 407 961 454
rect 878 401 973 407
rect 128 393 222 399
rect 128 327 140 393
rect 210 327 222 393
rect 128 321 222 327
rect 878 330 890 401
rect 961 330 973 401
rect 878 324 973 330
rect 1054 -158 1129 608
rect 1054 -221 1060 -158
rect 1123 -221 1129 -158
rect 1054 -233 1129 -221
use CNRATR_NCH_12C1F2  CNRATR_NCH_12C1F2_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 694 -1 0 2156
box -184 -124 2296 613
use CNRATR_NCH_12C1F2  CNRATR_NCH_12C1F2_1
timestamp 1695852000
transform 0 1 -56 -1 0 2156
box -184 -124 2296 613
<< labels >>
flabel locali 390 2310 470 2350 0 FreeSans 800 0 0 0 VDD
port 2 nsew
flabel locali 260 -240 390 -200 0 FreeSans 800 0 0 0 VSS
port 3 nsew
<< end >>
