*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/OTA_lpe.spi
#else
.include ../../../work/xsch/OTA.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  dc 1.8

VIN VIN VSS dc 0.9
V_DIFF VP VN ac 1



*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------

.save all

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 1 1 1 100p 20u 0


*tran 1n 20u 1n
ac dec 50 100 10G
settype decibel VO
plot vdb(VO) xlimit 1 100k ylabel 'small signal gain'
settype phase VO
plot cph(VO) xlimit 1 100k ylabel 'phase (in rad)'
let outd = 180/PI*cph(VO)
settype phase outd
plot outd xlimit 1 100k ylabel 'phase'

set gnuplot_terminal=png/quit
gnuplot {cicname}_loop_gain VO
gnuplot {cicname}_loop_phase outd

write


.endc

.end
