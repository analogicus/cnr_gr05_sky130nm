magic
tech sky130B
magscale 1 2
timestamp 1713514263
<< locali >>
rect 2202 8446 7660 8822
rect 4900 6221 4998 6230
rect 4900 6135 4912 6221
rect 4900 6132 4998 6135
rect 2946 -1422 3032 89
rect 6851 -1420 6937 89
rect 2944 -2160 4476 -1964
rect 5400 -2156 6940 -1966
rect 790 -10124 9086 -9978
<< viali >>
rect 4912 6135 4998 6221
rect 1977 4357 2155 4535
rect 7681 4369 7859 4547
rect 3118 -260 3308 -70
rect 6576 -260 6766 -70
<< metal1 >>
rect 4906 6227 5004 6233
rect 4900 6129 4906 6227
rect 5004 6129 5010 6227
rect 4906 6123 5004 6129
rect 7675 4547 7865 4559
rect 1971 4535 2161 4547
rect 1971 4357 1977 4535
rect 2155 4357 2161 4535
rect 1971 -70 2161 4357
rect 7675 4369 7681 4547
rect 7859 4369 7865 4547
rect 3112 -70 3314 -58
rect 1971 -260 3118 -70
rect 3308 -260 3314 -70
rect 3112 -272 3314 -260
rect 6570 -70 6772 -58
rect 7675 -70 7865 4369
rect 6570 -260 6576 -70
rect 6766 -260 7865 -70
rect 6570 -272 6772 -260
rect 4906 -1556 5004 -1550
rect 4896 -1654 4906 -1558
rect 4906 -1660 5004 -1654
<< via1 >>
rect 4906 6221 5004 6227
rect 4906 6135 4912 6221
rect 4912 6135 4998 6221
rect 4998 6135 5004 6221
rect 4906 6129 5004 6135
rect 4906 -1654 5004 -1556
<< metal2 >>
rect 4911 6227 4999 6231
rect 4900 6129 4906 6227
rect 5004 6129 5010 6227
rect 4911 6125 4999 6129
rect 4906 -1556 5004 -1547
rect 4900 -1654 4906 -1556
rect 5004 -1654 5010 -1556
rect 4906 -1663 5004 -1654
<< via2 >>
rect 4911 6134 4999 6222
rect 4906 -1654 5004 -1556
<< metal3 >>
rect 4906 6222 5004 6227
rect 4906 6134 4911 6222
rect 4999 6134 5004 6222
rect 4906 -1551 5004 6134
rect 4901 -1556 5009 -1551
rect 4901 -1654 4906 -1556
rect 5004 -1654 5009 -1556
rect 4901 -1659 5009 -1654
use IREF  IREF_0
timestamp 1713513383
transform 1 0 3800 0 1 -1114
box -3026 -8906 5302 1046
use PTAT  PTAT_0
timestamp 1713511997
transform 1 0 4270 0 1 180
box -4270 -180 5596 8590
<< labels >>
flabel locali 4604 8786 4754 8804 0 FreeSans 1600 0 0 0 VDD_1V8
port 3 nsew
flabel locali 7766 -10108 7968 -10042 0 FreeSans 1600 0 0 0 VSS
port 5 nsew
<< end >>
