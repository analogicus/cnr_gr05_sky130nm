magic
tech sky130B
timestamp 1713000619
<< nwell >>
rect -1100 -18 -1058 -13
<< pwell >>
rect -581 -1450 562 -1331
<< locali >>
rect -1099 709 1051 740
rect -1099 673 -48 709
rect -12 673 1051 709
rect -1099 636 1051 673
rect -1099 632 -1058 636
rect -1100 -18 -1058 632
rect -549 280 -518 283
rect 1001 -18 1051 636
rect -582 -790 -534 -109
rect 516 -122 562 -109
rect -581 -1331 -534 -790
rect 515 -1331 562 -122
rect -581 -1387 562 -1331
rect -581 -1413 -20 -1387
rect 6 -1413 562 -1387
rect -581 -1450 562 -1413
<< viali >>
rect -48 673 -12 709
rect -452 433 -426 459
rect 409 430 437 457
rect -84 294 -48 330
rect -1 297 29 327
rect -552 244 -516 280
rect 464 248 494 278
rect -455 -333 -423 -301
rect -26 -497 10 -461
rect -25 -589 7 -557
rect 407 -909 439 -877
rect -22 -1072 4 -1046
rect -23 -1165 9 -1133
rect -20 -1413 6 -1387
<< metal1 >>
rect -54 709 -6 712
rect -54 673 -48 709
rect -12 673 -6 709
rect -54 670 -6 673
rect -455 462 -423 465
rect -455 427 -423 430
rect -48 333 -12 670
rect 406 460 440 463
rect 406 424 440 427
rect -90 330 -12 333
rect -90 294 -84 330
rect -48 327 35 330
rect -48 297 -1 327
rect 29 297 35 327
rect -48 294 35 297
rect -90 291 -42 294
rect -558 280 -510 283
rect -558 244 -552 280
rect -516 244 -510 280
rect -558 241 -510 244
rect 461 278 497 284
rect 461 248 464 278
rect 494 248 497 278
rect -552 146 -516 241
rect -26 146 10 147
rect 461 146 497 248
rect -552 110 497 146
rect -458 -298 -420 -295
rect -461 -330 -458 -298
rect -420 -330 -417 -298
rect -461 -333 -455 -330
rect -423 -333 -417 -330
rect -461 -336 -417 -333
rect -26 -458 10 110
rect -32 -461 16 -458
rect -32 -497 -26 -461
rect 10 -497 16 -461
rect -32 -500 16 -497
rect -31 -557 13 -554
rect -31 -589 -25 -557
rect 7 -589 13 -557
rect -31 -592 13 -589
rect -25 -1046 7 -592
rect 401 -877 445 -874
rect 401 -880 407 -877
rect 439 -880 445 -877
rect 401 -912 404 -880
rect 442 -912 445 -880
rect 404 -915 442 -912
rect -25 -1072 -22 -1046
rect 4 -1072 7 -1046
rect -25 -1078 7 -1072
rect -29 -1133 15 -1130
rect -29 -1165 -23 -1133
rect 9 -1165 15 -1133
rect -29 -1168 15 -1165
rect -23 -1387 9 -1168
rect -23 -1413 -20 -1387
rect 6 -1413 9 -1387
rect -23 -1419 9 -1413
<< via1 >>
rect -455 459 -423 462
rect -455 433 -452 459
rect -452 433 -426 459
rect -426 433 -423 459
rect -455 430 -423 433
rect 406 457 440 460
rect 406 430 409 457
rect 409 430 437 457
rect 437 430 440 457
rect 406 427 440 430
rect -458 -301 -420 -298
rect -458 -330 -455 -301
rect -455 -330 -423 -301
rect -423 -330 -420 -301
rect 404 -909 407 -880
rect 407 -909 439 -880
rect 439 -909 442 -880
rect 404 -912 442 -909
<< metal2 >>
rect -458 430 -455 462
rect -423 430 -420 462
rect -455 -298 -423 430
rect 403 427 406 460
rect 440 427 443 460
rect -461 -330 -458 -298
rect -420 -330 -417 -298
rect 406 -880 440 427
rect 401 -912 404 -880
rect 442 -912 445 -880
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 -1 502 1 0 -1309
box -92 -62 668 1084
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_1
timestamp 1695852000
transform 0 -1 502 1 0 -733
box -92 -62 668 1084
use CNRATR_PCH_2C12F0  CNRATR_PCH_2C12F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 -1 -23 1 0 30
box -92 -62 668 1084
use CNRATR_PCH_2C12F0  CNRATR_PCH_2C12F0_1
timestamp 1695852000
transform 0 -1 992 1 0 30
box -92 -62 668 1084
<< labels >>
flabel locali 106 677 180 712 0 FreeSans 800 0 0 0 VDD_1V8
port 1 nsew
flabel locali 159 -1434 233 -1399 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel metal1 -24 -283 2 -257 0 FreeSans 200 0 0 0 O
port 4 nsew
flabel metal2 -450 -91 -424 -65 0 FreeSans 200 0 0 0 A
port 3 nsew
flabel metal2 407 -104 433 -78 0 FreeSans 200 0 0 0 B
port 5 nsew
<< end >>
