magic
tech sky130B
magscale 1 2
timestamp 1713000619
<< nwell >>
rect -2200 -36 -2116 -26
<< pwell >>
rect -1162 -2900 1124 -2662
<< locali >>
rect -2198 1418 2102 1480
rect -2198 1346 -96 1418
rect -24 1346 2102 1418
rect -2198 1272 2102 1346
rect -2198 1264 -2116 1272
rect -2200 -36 -2116 1264
rect -1098 560 -1036 566
rect 2002 -36 2102 1272
rect -1164 -1580 -1068 -218
rect 1032 -244 1124 -218
rect -1162 -2662 -1068 -1580
rect 1030 -2662 1124 -244
rect -1162 -2774 1124 -2662
rect -1162 -2826 -40 -2774
rect 12 -2826 1124 -2774
rect -1162 -2900 1124 -2826
<< viali >>
rect -96 1346 -24 1418
rect -904 866 -852 918
rect 819 860 874 915
rect -168 588 -96 660
rect -2 594 58 654
rect -1104 488 -1032 560
rect 928 496 988 556
rect -910 -666 -846 -602
rect -52 -994 20 -922
rect -50 -1178 14 -1114
rect 814 -1818 878 -1754
rect -44 -2144 8 -2092
rect -46 -2330 18 -2266
rect -40 -2826 12 -2774
<< metal1 >>
rect -108 1418 -12 1424
rect -108 1346 -96 1418
rect -24 1346 -12 1418
rect -108 1340 -12 1346
rect -910 924 -846 930
rect -910 854 -846 860
rect -96 666 -24 1340
rect 813 921 880 927
rect 813 848 880 854
rect -180 660 -24 666
rect -180 588 -168 660
rect -96 654 70 660
rect -96 594 -2 654
rect 58 594 70 654
rect -96 588 70 594
rect -180 582 -84 588
rect -1116 560 -1020 566
rect -1116 488 -1104 560
rect -1032 488 -1020 560
rect -1116 482 -1020 488
rect 922 556 994 568
rect 922 496 928 556
rect 988 496 994 556
rect -1104 292 -1032 482
rect -52 292 20 294
rect 922 292 994 496
rect -1104 220 994 292
rect -916 -596 -840 -590
rect -922 -660 -916 -596
rect -840 -660 -834 -596
rect -922 -666 -910 -660
rect -846 -666 -834 -660
rect -922 -672 -834 -666
rect -52 -916 20 220
rect -64 -922 32 -916
rect -64 -994 -52 -922
rect 20 -994 32 -922
rect -64 -1000 32 -994
rect -62 -1114 26 -1108
rect -62 -1178 -50 -1114
rect 14 -1178 26 -1114
rect -62 -1184 26 -1178
rect -50 -2092 14 -1184
rect 802 -1754 890 -1748
rect 802 -1760 814 -1754
rect 878 -1760 890 -1754
rect 802 -1824 808 -1760
rect 884 -1824 890 -1760
rect 808 -1830 884 -1824
rect -50 -2144 -44 -2092
rect 8 -2144 14 -2092
rect -50 -2156 14 -2144
rect -58 -2266 30 -2260
rect -58 -2330 -46 -2266
rect 18 -2330 30 -2266
rect -58 -2336 30 -2330
rect -46 -2774 18 -2336
rect -46 -2826 -40 -2774
rect 12 -2826 18 -2774
rect -46 -2838 18 -2826
<< via1 >>
rect -910 918 -846 924
rect -910 866 -904 918
rect -904 866 -852 918
rect -852 866 -846 918
rect -910 860 -846 866
rect 813 915 880 921
rect 813 860 819 915
rect 819 860 874 915
rect 874 860 880 915
rect 813 854 880 860
rect -916 -602 -840 -596
rect -916 -660 -910 -602
rect -910 -660 -846 -602
rect -846 -660 -840 -602
rect 808 -1818 814 -1760
rect 814 -1818 878 -1760
rect 878 -1818 884 -1760
rect 808 -1824 884 -1818
<< metal2 >>
rect -916 860 -910 924
rect -846 860 -840 924
rect -910 -596 -846 860
rect 807 854 813 921
rect 880 854 886 921
rect -922 -660 -916 -596
rect -840 -660 -834 -596
rect 813 -1760 880 854
rect 802 -1824 808 -1760
rect 884 -1824 890 -1760
rect 813 -1825 880 -1824
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 -1 1004 1 0 -2618
box -184 -124 1336 2168
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_1
timestamp 1695852000
transform 0 -1 1004 1 0 -1466
box -184 -124 1336 2168
use CNRATR_PCH_2C12F0  CNRATR_PCH_2C12F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 -1 -46 1 0 60
box -184 -124 1336 2168
use CNRATR_PCH_2C12F0  CNRATR_PCH_2C12F0_1
timestamp 1695852000
transform 0 -1 1984 1 0 60
box -184 -124 1336 2168
<< labels >>
flabel locali 212 1354 360 1424 0 FreeSans 1600 0 0 0 VDD_1V8
port 1 nsew
flabel locali 318 -2868 466 -2798 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 -48 -566 4 -514 0 FreeSans 400 0 0 0 O
port 4 nsew
flabel metal2 -900 -182 -848 -130 0 FreeSans 400 0 0 0 A
port 3 nsew
flabel metal2 814 -208 866 -156 0 FreeSans 400 0 0 0 B
port 5 nsew
<< end >>
