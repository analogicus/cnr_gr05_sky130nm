*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_05_lpe.spi
#else
.include ../../../work/xsch/CNR_GR05.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0 dc 0
VDD_1V8  VDD_1V8  0 dc 1.8
*VP VP 0 dc 1.2

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VP VN VSS VDD_1V8 CNR_GR05


*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
*.save ${VPORTS}
#endif
.save all
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 1 1 1 100p 2n 0

#ifdef Debug
tran 10p 1n 1p
*quit
#else
tran 10p 100n 1p
write
quit
#endif

.endc

.end