magic
tech sky130B
timestamp 1713355520
<< locali >>
rect 2118 2269 2790 2299
rect 350 1994 401 1995
rect 350 1898 459 1994
rect 1497 1898 2198 1994
rect 350 1418 401 1898
rect 350 1322 461 1418
rect 350 842 401 1322
rect 350 746 458 842
rect 2018 558 2133 654
rect 2016 -117 2212 78
<< viali >>
rect 978 1935 1004 1961
rect 975 1770 1007 1802
rect 974 1647 1000 1673
rect 535 1514 567 1546
rect 971 1194 1003 1226
rect 974 1078 1000 1104
rect 1403 938 1435 970
rect 538 433 564 459
rect 1406 434 1432 460
rect 463 271 495 305
rect 1483 275 1509 301
rect 471 174 503 206
rect 1478 174 1510 206
rect 474 17 500 43
rect 1481 17 1507 43
<< metal1 >>
rect 975 1961 1007 1967
rect 975 1935 978 1961
rect 1004 1935 1007 1961
rect 975 1805 1007 1935
rect 969 1802 1013 1805
rect 969 1770 975 1802
rect 1007 1770 1013 1802
rect 969 1767 1013 1770
rect 971 1673 1003 1679
rect 971 1647 974 1673
rect 1000 1647 1003 1673
rect 529 1546 573 1549
rect 529 1514 535 1546
rect 567 1514 573 1546
rect 529 1511 573 1514
rect 535 733 567 1511
rect 971 1229 1003 1647
rect 965 1226 1009 1229
rect 965 1194 971 1226
rect 1003 1194 1009 1226
rect 965 1191 1009 1194
rect 971 1104 1003 1110
rect 971 1078 974 1104
rect 1000 1078 1003 1104
rect 971 900 1003 1078
rect 2390 1010 2438 1137
rect 2567 1095 2599 1098
rect 2567 1060 2599 1063
rect 1397 970 1441 973
rect 1397 938 1403 970
rect 1435 938 1441 970
rect 1397 935 1441 938
rect 968 868 971 900
rect 1003 868 1006 900
rect 535 670 613 733
rect 535 462 567 670
rect 532 459 570 462
rect 532 433 538 459
rect 564 433 570 459
rect 532 430 570 433
rect 460 305 498 311
rect 460 271 463 305
rect 495 304 498 305
rect 971 304 1003 868
rect 1403 736 1435 935
rect 1403 666 1493 736
rect 1403 460 1435 666
rect 1403 434 1406 460
rect 1432 434 1435 460
rect 1403 428 1435 434
rect 495 301 1515 304
rect 495 275 1483 301
rect 1509 275 1515 301
rect 495 272 1515 275
rect 495 271 498 272
rect 460 265 498 271
rect 465 206 509 209
rect 465 174 471 206
rect 503 174 509 206
rect 465 171 509 174
rect 1472 206 1516 209
rect 1472 174 1478 206
rect 1510 174 1516 206
rect 1472 171 1516 174
rect 471 43 503 171
rect 471 17 474 43
rect 500 17 503 43
rect 471 11 503 17
rect 1478 43 1510 171
rect 1478 17 1481 43
rect 1507 17 1510 43
rect 1478 11 1510 17
<< via1 >>
rect 2567 1063 2599 1095
rect 971 868 1003 900
<< metal2 >>
rect 1990 1063 2567 1095
rect 2599 1063 2602 1095
rect 971 900 1003 903
rect 1990 900 2022 1063
rect 1003 868 2022 900
rect 971 865 1003 868
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 -1 2007 1 0 30
box -92 -62 668 1084
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_1
timestamp 1695852000
transform 0 -1 992 1 0 30
box -92 -62 668 1084
use CNRATR_PCH_2C12F0  CNRATR_PCH_2C12F0_0 ~/aicex/ip/cnr_gr05_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 474 -1 0 1946
box -92 -62 668 1084
use CNRATR_PCH_2C12F0  CNRATR_PCH_2C12F0_1
timestamp 1695852000
transform 0 1 474 -1 0 1370
box -92 -62 668 1084
use INV  INV_0
timestamp 1712998694
transform 1 0 2164 0 1 2
box -92 -119 670 2277
<< labels >>
flabel locali 2423 2286 2448 2293 0 FreeSans 200 0 0 0 VDD_1V8
port 1 nsew
flabel locali 2044 -81 2077 -41 0 FreeSans 200 0 0 0 VSS
port 2 nsew
flabel metal1 2400 1106 2416 1123 0 FreeSans 200 0 0 0 O
port 4 nsew
flabel metal1 1450 683 1472 717 0 FreeSans 200 0 0 0 B
port 5 nsew
flabel metal1 579 686 600 713 0 FreeSans 200 0 0 0 A
port 3 nsew
<< end >>
